module NOT_Gate(input in,
				output out );

    assign out = ~in;
    
endmodule
